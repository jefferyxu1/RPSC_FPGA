module card1();

endmodule